// Module to control branch operations

module branch_control(BranchOp,zero,pc_in,pc_out);
    
endmodule