module and_module(a,b,result); // AND gate
    output [7:0] result;
    
    assign result = a & b; // bitwise AND
endmodule