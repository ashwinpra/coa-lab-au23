// Module to control stack operations

module stack_control(StackOp);
    input [2:0] StackOp;

    
endmodule