// arithmetic right shift 
module a_rshift(A, Q, Q_1, out); 
    input [7:0] A, Q;
    input Q_1; 
    output [7:0] out;
endmodule