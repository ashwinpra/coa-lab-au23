module move (a,result); // move module
    input [7:0] a;
    output [7:0] result;
    
    assign result = a; // move a to result
endmodule